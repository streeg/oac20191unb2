DecoderIP_inst : DecoderIP PORT MAP (
		data	 => data_sig
	);
