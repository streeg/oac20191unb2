comparador_inst : comparador PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		aeb	 => aeb_sig
	);
